//Controller

/*
module controller(
						input wire [5:0] opcode,
						output reg regfile,
						output reg alucunt,
						output reg alusrc,
						output reg memwrite,
						output reg memread,
						output reg memtoreg,
						output reg pcsrc,
						output reg regdist);
						
						
//Send one 8 bit output reg through the pipeline, each bit representing a different control bit. 
*/