//Test to blink LED

module blink(LEDG);

	output[7:0] LEDG;
	
	assign LEDG[0] = 1'b0;
	
endmodule


	