library verilog;
use verilog.vl_types.all;
entity registerfile_vlg_vec_tst is
end registerfile_vlg_vec_tst;
