library verilog;
use verilog.vl_types.all;
entity simpleregister_vlg_vec_tst is
end simpleregister_vlg_vec_tst;
